library IEEE;
use IEEE.STD_LOGIC_1164.all;

library IEEE_PROPOSED;
use IEEE_PROPOSED.FIXED_PKG.ALL;

package Trigo is
	function sin (val: INTEGER) return sfixed is
		variable ret : sfixed(11 downto -20);
	begin
		case val is
			when 0 =>
				ret := to_sfixed(0.0, ret);
			when 1 =>
				ret := to_sfixed(0.01745241, ret);
			when 2 =>
				ret := to_sfixed(0.0348995, ret);
			when 3 =>
				ret := to_sfixed(0.05233596, ret);
			when 4 =>
				ret := to_sfixed(0.06975647, ret);
			when 5 =>
				ret := to_sfixed(0.08715574, ret);
			when 6 =>
				ret := to_sfixed(0.10452846, ret);
			when 7 =>
				ret := to_sfixed(0.12186934, ret);
			when 8 =>
				ret := to_sfixed(0.1391731, ret);
			when 9 =>
				ret := to_sfixed(0.15643447, ret);
			when 10 =>
				ret := to_sfixed(0.17364818, ret);
			when 11 =>
				ret := to_sfixed(0.190809, ret);
			when 12 =>
				ret := to_sfixed(0.20791169, ret);
			when 13 =>
				ret := to_sfixed(0.22495105, ret);
			when 14 =>
				ret := to_sfixed(0.2419219, ret);
			when 15 =>
				ret := to_sfixed(0.25881905, ret);
			when 16 =>
				ret := to_sfixed(0.27563736, ret);
			when 17 =>
				ret := to_sfixed(0.2923717, ret);
			when 18 =>
				ret := to_sfixed(0.30901699, ret);
			when 19 =>
				ret := to_sfixed(0.32556815, ret);
			when 20 =>
				ret := to_sfixed(0.34202014, ret);
			when 21 =>
				ret := to_sfixed(0.35836795, ret);
			when 22 =>
				ret := to_sfixed(0.37460659, ret);
			when 23 =>
				ret := to_sfixed(0.39073113, ret);
			when 24 =>
				ret := to_sfixed(0.40673664, ret);
			when 25 =>
				ret := to_sfixed(0.42261826, ret);
			when 26 =>
				ret := to_sfixed(0.43837115, ret);
			when 27 =>
				ret := to_sfixed(0.4539905, ret);
			when 28 =>
				ret := to_sfixed(0.46947156, ret);
			when 29 =>
				ret := to_sfixed(0.48480962, ret);
			when 30 =>
				ret := to_sfixed(0.5, ret);
			when 31 =>
				ret := to_sfixed(0.51503807, ret);
			when 32 =>
				ret := to_sfixed(0.52991926, ret);
			when 33 =>
				ret := to_sfixed(0.54463904, ret);
			when 34 =>
				ret := to_sfixed(0.5591929, ret);
			when 35 =>
				ret := to_sfixed(0.57357644, ret);
			when 36 =>
				ret := to_sfixed(0.58778525, ret);
			when 37 =>
				ret := to_sfixed(0.60181502, ret);
			when 38 =>
				ret := to_sfixed(0.61566148, ret);
			when 39 =>
				ret := to_sfixed(0.62932039, ret);
			when 40 =>
				ret := to_sfixed(0.64278761, ret);
			when 41 =>
				ret := to_sfixed(0.65605903, ret);
			when 42 =>
				ret := to_sfixed(0.66913061, ret);
			when 43 =>
				ret := to_sfixed(0.68199836, ret);
			when 44 =>
				ret := to_sfixed(0.69465837, ret);
			when 45 =>
				ret := to_sfixed(0.70710678, ret);
			when 46 =>
				ret := to_sfixed(0.7193398, ret);
			when 47 =>
				ret := to_sfixed(0.7313537, ret);
			when 48 =>
				ret := to_sfixed(0.74314483, ret);
			when 49 =>
				ret := to_sfixed(0.75470958, ret);
			when 50 =>
				ret := to_sfixed(0.76604444, ret);
			when 51 =>
				ret := to_sfixed(0.77714596, ret);
			when 52 =>
				ret := to_sfixed(0.78801075, ret);
			when 53 =>
				ret := to_sfixed(0.79863551, ret);
			when 54 =>
				ret := to_sfixed(0.80901699, ret);
			when 55 =>
				ret := to_sfixed(0.81915204, ret);
			when 56 =>
				ret := to_sfixed(0.82903757, ret);
			when 57 =>
				ret := to_sfixed(0.83867057, ret);
			when 58 =>
				ret := to_sfixed(0.8480481, ret);
			when 59 =>
				ret := to_sfixed(0.8571673, ret);
			when 60 =>
				ret := to_sfixed(0.8660254, ret);
			when 61 =>
				ret := to_sfixed(0.87461971, ret);
			when 62 =>
				ret := to_sfixed(0.88294759, ret);
			when 63 =>
				ret := to_sfixed(0.89100652, ret);
			when 64 =>
				ret := to_sfixed(0.89879405, ret);
			when 65 =>
				ret := to_sfixed(0.90630779, ret);
			when 66 =>
				ret := to_sfixed(0.91354546, ret);
			when 67 =>
				ret := to_sfixed(0.92050485, ret);
			when 68 =>
				ret := to_sfixed(0.92718385, ret);
			when 69 =>
				ret := to_sfixed(0.93358043, ret);
			when 70 =>
				ret := to_sfixed(0.93969262, ret);
			when 71 =>
				ret := to_sfixed(0.94551858, ret);
			when 72 =>
				ret := to_sfixed(0.95105652, ret);
			when 73 =>
				ret := to_sfixed(0.95630476, ret);
			when 74 =>
				ret := to_sfixed(0.9612617, ret);
			when 75 =>
				ret := to_sfixed(0.96592583, ret);
			when 76 =>
				ret := to_sfixed(0.97029573, ret);
			when 77 =>
				ret := to_sfixed(0.97437006, ret);
			when 78 =>
				ret := to_sfixed(0.9781476, ret);
			when 79 =>
				ret := to_sfixed(0.98162718, ret);
			when 80 =>
				ret := to_sfixed(0.98480775, ret);
			when 81 =>
				ret := to_sfixed(0.98768834, ret);
			when 82 =>
				ret := to_sfixed(0.99026807, ret);
			when 83 =>
				ret := to_sfixed(0.99254615, ret);
			when 84 =>
				ret := to_sfixed(0.9945219, ret);
			when 85 =>
				ret := to_sfixed(0.9961947, ret);
			when 86 =>
				ret := to_sfixed(0.99756405, ret);
			when 87 =>
				ret := to_sfixed(0.99862953, ret);
			when 88 =>
				ret := to_sfixed(0.99939083, ret);
			when 89 =>
				ret := to_sfixed(0.9998477, ret);
			when 90 =>
				ret := to_sfixed(1.0, ret);
			when 91 =>
				ret := to_sfixed(0.9998477, ret);
			when 92 =>
				ret := to_sfixed(0.99939083, ret);
			when 93 =>
				ret := to_sfixed(0.99862953, ret);
			when 94 =>
				ret := to_sfixed(0.99756405, ret);
			when 95 =>
				ret := to_sfixed(0.9961947, ret);
			when 96 =>
				ret := to_sfixed(0.9945219, ret);
			when 97 =>
				ret := to_sfixed(0.99254615, ret);
			when 98 =>
				ret := to_sfixed(0.99026807, ret);
			when 99 =>
				ret := to_sfixed(0.98768834, ret);
			when 100 =>
				ret := to_sfixed(0.98480775, ret);
			when 101 =>
				ret := to_sfixed(0.98162718, ret);
			when 102 =>
				ret := to_sfixed(0.9781476, ret);
			when 103 =>
				ret := to_sfixed(0.97437006, ret);
			when 104 =>
				ret := to_sfixed(0.97029573, ret);
			when 105 =>
				ret := to_sfixed(0.96592583, ret);
			when 106 =>
				ret := to_sfixed(0.9612617, ret);
			when 107 =>
				ret := to_sfixed(0.95630476, ret);
			when 108 =>
				ret := to_sfixed(0.95105652, ret);
			when 109 =>
				ret := to_sfixed(0.94551858, ret);
			when 110 =>
				ret := to_sfixed(0.93969262, ret);
			when 111 =>
				ret := to_sfixed(0.93358043, ret);
			when 112 =>
				ret := to_sfixed(0.92718385, ret);
			when 113 =>
				ret := to_sfixed(0.92050485, ret);
			when 114 =>
				ret := to_sfixed(0.91354546, ret);
			when 115 =>
				ret := to_sfixed(0.90630779, ret);
			when 116 =>
				ret := to_sfixed(0.89879405, ret);
			when 117 =>
				ret := to_sfixed(0.89100652, ret);
			when 118 =>
				ret := to_sfixed(0.88294759, ret);
			when 119 =>
				ret := to_sfixed(0.87461971, ret);
			when 120 =>
				ret := to_sfixed(0.8660254, ret);
			when 121 =>
				ret := to_sfixed(0.8571673, ret);
			when 122 =>
				ret := to_sfixed(0.8480481, ret);
			when 123 =>
				ret := to_sfixed(0.83867057, ret);
			when 124 =>
				ret := to_sfixed(0.82903757, ret);
			when 125 =>
				ret := to_sfixed(0.81915204, ret);
			when 126 =>
				ret := to_sfixed(0.80901699, ret);
			when 127 =>
				ret := to_sfixed(0.79863551, ret);
			when 128 =>
				ret := to_sfixed(0.78801075, ret);
			when 129 =>
				ret := to_sfixed(0.77714596, ret);
			when 130 =>
				ret := to_sfixed(0.76604444, ret);
			when 131 =>
				ret := to_sfixed(0.75470958, ret);
			when 132 =>
				ret := to_sfixed(0.74314483, ret);
			when 133 =>
				ret := to_sfixed(0.7313537, ret);
			when 134 =>
				ret := to_sfixed(0.7193398, ret);
			when 135 =>
				ret := to_sfixed(0.70710678, ret);
			when 136 =>
				ret := to_sfixed(0.69465837, ret);
			when 137 =>
				ret := to_sfixed(0.68199836, ret);
			when 138 =>
				ret := to_sfixed(0.66913061, ret);
			when 139 =>
				ret := to_sfixed(0.65605903, ret);
			when 140 =>
				ret := to_sfixed(0.64278761, ret);
			when 141 =>
				ret := to_sfixed(0.62932039, ret);
			when 142 =>
				ret := to_sfixed(0.61566148, ret);
			when 143 =>
				ret := to_sfixed(0.60181502, ret);
			when 144 =>
				ret := to_sfixed(0.58778525, ret);
			when 145 =>
				ret := to_sfixed(0.57357644, ret);
			when 146 =>
				ret := to_sfixed(0.5591929, ret);
			when 147 =>
				ret := to_sfixed(0.54463904, ret);
			when 148 =>
				ret := to_sfixed(0.52991926, ret);
			when 149 =>
				ret := to_sfixed(0.51503807, ret);
			when 150 =>
				ret := to_sfixed(0.5, ret);
			when 151 =>
				ret := to_sfixed(0.48480962, ret);
			when 152 =>
				ret := to_sfixed(0.46947156, ret);
			when 153 =>
				ret := to_sfixed(0.4539905, ret);
			when 154 =>
				ret := to_sfixed(0.43837115, ret);
			when 155 =>
				ret := to_sfixed(0.42261826, ret);
			when 156 =>
				ret := to_sfixed(0.40673664, ret);
			when 157 =>
				ret := to_sfixed(0.39073113, ret);
			when 158 =>
				ret := to_sfixed(0.37460659, ret);
			when 159 =>
				ret := to_sfixed(0.35836795, ret);
			when 160 =>
				ret := to_sfixed(0.34202014, ret);
			when 161 =>
				ret := to_sfixed(0.32556815, ret);
			when 162 =>
				ret := to_sfixed(0.30901699, ret);
			when 163 =>
				ret := to_sfixed(0.2923717, ret);
			when 164 =>
				ret := to_sfixed(0.27563736, ret);
			when 165 =>
				ret := to_sfixed(0.25881905, ret);
			when 166 =>
				ret := to_sfixed(0.2419219, ret);
			when 167 =>
				ret := to_sfixed(0.22495105, ret);
			when 168 =>
				ret := to_sfixed(0.20791169, ret);
			when 169 =>
				ret := to_sfixed(0.190809, ret);
			when 170 =>
				ret := to_sfixed(0.17364818, ret);
			when 171 =>
				ret := to_sfixed(0.15643447, ret);
			when 172 =>
				ret := to_sfixed(0.1391731, ret);
			when 173 =>
				ret := to_sfixed(0.12186934, ret);
			when 174 =>
				ret := to_sfixed(0.10452846, ret);
			when 175 =>
				ret := to_sfixed(0.08715574, ret);
			when 176 =>
				ret := to_sfixed(0.06975647, ret);
			when 177 =>
				ret := to_sfixed(0.05233596, ret);
			when 178 =>
				ret := to_sfixed(0.0348995, ret);
			when 179 =>
				ret := to_sfixed(0.01745241, ret);
			when others =>
				ret := to_sfixed(0.0, ret);
		end case;
		return ret; 
	end sin;

	function cos (val: INTEGER) return sfixed is
		variable ret : sfixed(11 downto -20);
	begin
		case val is
			when 0 =>
				ret := to_sfixed(1.0, ret);
			when 1 =>
				ret := to_sfixed(0.9998477, ret);
			when 2 =>
				ret := to_sfixed(0.99939083, ret);
			when 3 =>
				ret := to_sfixed(0.99862953, ret);
			when 4 =>
				ret := to_sfixed(0.99756405, ret);
			when 5 =>
				ret := to_sfixed(0.9961947, ret);
			when 6 =>
				ret := to_sfixed(0.9945219, ret);
			when 7 =>
				ret := to_sfixed(0.99254615, ret);
			when 8 =>
				ret := to_sfixed(0.99026807, ret);
			when 9 =>
				ret := to_sfixed(0.98768834, ret);
			when 10 =>
				ret := to_sfixed(0.98480775, ret);
			when 11 =>
				ret := to_sfixed(0.98162718, ret);
			when 12 =>
				ret := to_sfixed(0.9781476, ret);
			when 13 =>
				ret := to_sfixed(0.97437006, ret);
			when 14 =>
				ret := to_sfixed(0.97029573, ret);
			when 15 =>
				ret := to_sfixed(0.96592583, ret);
			when 16 =>
				ret := to_sfixed(0.9612617, ret);
			when 17 =>
				ret := to_sfixed(0.95630476, ret);
			when 18 =>
				ret := to_sfixed(0.95105652, ret);
			when 19 =>
				ret := to_sfixed(0.94551858, ret);
			when 20 =>
				ret := to_sfixed(0.93969262, ret);
			when 21 =>
				ret := to_sfixed(0.93358043, ret);
			when 22 =>
				ret := to_sfixed(0.92718385, ret);
			when 23 =>
				ret := to_sfixed(0.92050485, ret);
			when 24 =>
				ret := to_sfixed(0.91354546, ret);
			when 25 =>
				ret := to_sfixed(0.90630779, ret);
			when 26 =>
				ret := to_sfixed(0.89879405, ret);
			when 27 =>
				ret := to_sfixed(0.89100652, ret);
			when 28 =>
				ret := to_sfixed(0.88294759, ret);
			when 29 =>
				ret := to_sfixed(0.87461971, ret);
			when 30 =>
				ret := to_sfixed(0.8660254, ret);
			when 31 =>
				ret := to_sfixed(0.8571673, ret);
			when 32 =>
				ret := to_sfixed(0.8480481, ret);
			when 33 =>
				ret := to_sfixed(0.83867057, ret);
			when 34 =>
				ret := to_sfixed(0.82903757, ret);
			when 35 =>
				ret := to_sfixed(0.81915204, ret);
			when 36 =>
				ret := to_sfixed(0.80901699, ret);
			when 37 =>
				ret := to_sfixed(0.79863551, ret);
			when 38 =>
				ret := to_sfixed(0.78801075, ret);
			when 39 =>
				ret := to_sfixed(0.77714596, ret);
			when 40 =>
				ret := to_sfixed(0.76604444, ret);
			when 41 =>
				ret := to_sfixed(0.75470958, ret);
			when 42 =>
				ret := to_sfixed(0.74314483, ret);
			when 43 =>
				ret := to_sfixed(0.7313537, ret);
			when 44 =>
				ret := to_sfixed(0.7193398, ret);
			when 45 =>
				ret := to_sfixed(0.70710678, ret);
			when 46 =>
				ret := to_sfixed(0.69465837, ret);
			when 47 =>
				ret := to_sfixed(0.68199836, ret);
			when 48 =>
				ret := to_sfixed(0.66913061, ret);
			when 49 =>
				ret := to_sfixed(0.65605903, ret);
			when 50 =>
				ret := to_sfixed(0.64278761, ret);
			when 51 =>
				ret := to_sfixed(0.62932039, ret);
			when 52 =>
				ret := to_sfixed(0.61566148, ret);
			when 53 =>
				ret := to_sfixed(0.60181502, ret);
			when 54 =>
				ret := to_sfixed(0.58778525, ret);
			when 55 =>
				ret := to_sfixed(0.57357644, ret);
			when 56 =>
				ret := to_sfixed(0.5591929, ret);
			when 57 =>
				ret := to_sfixed(0.54463904, ret);
			when 58 =>
				ret := to_sfixed(0.52991926, ret);
			when 59 =>
				ret := to_sfixed(0.51503807, ret);
			when 60 =>
				ret := to_sfixed(0.5, ret);
			when 61 =>
				ret := to_sfixed(0.48480962, ret);
			when 62 =>
				ret := to_sfixed(0.46947156, ret);
			when 63 =>
				ret := to_sfixed(0.4539905, ret);
			when 64 =>
				ret := to_sfixed(0.43837115, ret);
			when 65 =>
				ret := to_sfixed(0.42261826, ret);
			when 66 =>
				ret := to_sfixed(0.40673664, ret);
			when 67 =>
				ret := to_sfixed(0.39073113, ret);
			when 68 =>
				ret := to_sfixed(0.37460659, ret);
			when 69 =>
				ret := to_sfixed(0.35836795, ret);
			when 70 =>
				ret := to_sfixed(0.34202014, ret);
			when 71 =>
				ret := to_sfixed(0.32556815, ret);
			when 72 =>
				ret := to_sfixed(0.30901699, ret);
			when 73 =>
				ret := to_sfixed(0.2923717, ret);
			when 74 =>
				ret := to_sfixed(0.27563736, ret);
			when 75 =>
				ret := to_sfixed(0.25881905, ret);
			when 76 =>
				ret := to_sfixed(0.2419219, ret);
			when 77 =>
				ret := to_sfixed(0.22495105, ret);
			when 78 =>
				ret := to_sfixed(0.20791169, ret);
			when 79 =>
				ret := to_sfixed(0.190809, ret);
			when 80 =>
				ret := to_sfixed(0.17364818, ret);
			when 81 =>
				ret := to_sfixed(0.15643447, ret);
			when 82 =>
				ret := to_sfixed(0.1391731, ret);
			when 83 =>
				ret := to_sfixed(0.12186934, ret);
			when 84 =>
				ret := to_sfixed(0.10452846, ret);
			when 85 =>
				ret := to_sfixed(0.08715574, ret);
			when 86 =>
				ret := to_sfixed(0.06975647, ret);
			when 87 =>
				ret := to_sfixed(0.05233596, ret);
			when 88 =>
				ret := to_sfixed(0.0348995, ret);
			when 89 =>
				ret := to_sfixed(0.01745241, ret);
			when 90 =>
				ret := to_sfixed(0.0, ret);
			when 91 =>
				ret := to_sfixed(-0.01745241, ret);
			when 92 =>
				ret := to_sfixed(-0.0348995, ret);
			when 93 =>
				ret := to_sfixed(-0.05233596, ret);
			when 94 =>
				ret := to_sfixed(-0.06975647, ret);
			when 95 =>
				ret := to_sfixed(-0.08715574, ret);
			when 96 =>
				ret := to_sfixed(-0.10452846, ret);
			when 97 =>
				ret := to_sfixed(-0.12186934, ret);
			when 98 =>
				ret := to_sfixed(-0.1391731, ret);
			when 99 =>
				ret := to_sfixed(-0.15643447, ret);
			when 100 =>
				ret := to_sfixed(-0.17364818, ret);
			when 101 =>
				ret := to_sfixed(-0.190809, ret);
			when 102 =>
				ret := to_sfixed(-0.20791169, ret);
			when 103 =>
				ret := to_sfixed(-0.22495105, ret);
			when 104 =>
				ret := to_sfixed(-0.2419219, ret);
			when 105 =>
				ret := to_sfixed(-0.25881905, ret);
			when 106 =>
				ret := to_sfixed(-0.27563736, ret);
			when 107 =>
				ret := to_sfixed(-0.2923717, ret);
			when 108 =>
				ret := to_sfixed(-0.30901699, ret);
			when 109 =>
				ret := to_sfixed(-0.32556815, ret);
			when 110 =>
				ret := to_sfixed(-0.34202014, ret);
			when 111 =>
				ret := to_sfixed(-0.35836795, ret);
			when 112 =>
				ret := to_sfixed(-0.37460659, ret);
			when 113 =>
				ret := to_sfixed(-0.39073113, ret);
			when 114 =>
				ret := to_sfixed(-0.40673664, ret);
			when 115 =>
				ret := to_sfixed(-0.42261826, ret);
			when 116 =>
				ret := to_sfixed(-0.43837115, ret);
			when 117 =>
				ret := to_sfixed(-0.4539905, ret);
			when 118 =>
				ret := to_sfixed(-0.46947156, ret);
			when 119 =>
				ret := to_sfixed(-0.48480962, ret);
			when 120 =>
				ret := to_sfixed(-0.5, ret);
			when 121 =>
				ret := to_sfixed(-0.51503807, ret);
			when 122 =>
				ret := to_sfixed(-0.52991926, ret);
			when 123 =>
				ret := to_sfixed(-0.54463904, ret);
			when 124 =>
				ret := to_sfixed(-0.5591929, ret);
			when 125 =>
				ret := to_sfixed(-0.57357644, ret);
			when 126 =>
				ret := to_sfixed(-0.58778525, ret);
			when 127 =>
				ret := to_sfixed(-0.60181502, ret);
			when 128 =>
				ret := to_sfixed(-0.61566148, ret);
			when 129 =>
				ret := to_sfixed(-0.62932039, ret);
			when 130 =>
				ret := to_sfixed(-0.64278761, ret);
			when 131 =>
				ret := to_sfixed(-0.65605903, ret);
			when 132 =>
				ret := to_sfixed(-0.66913061, ret);
			when 133 =>
				ret := to_sfixed(-0.68199836, ret);
			when 134 =>
				ret := to_sfixed(-0.69465837, ret);
			when 135 =>
				ret := to_sfixed(-0.70710678, ret);
			when 136 =>
				ret := to_sfixed(-0.7193398, ret);
			when 137 =>
				ret := to_sfixed(-0.7313537, ret);
			when 138 =>
				ret := to_sfixed(-0.74314483, ret);
			when 139 =>
				ret := to_sfixed(-0.75470958, ret);
			when 140 =>
				ret := to_sfixed(-0.76604444, ret);
			when 141 =>
				ret := to_sfixed(-0.77714596, ret);
			when 142 =>
				ret := to_sfixed(-0.78801075, ret);
			when 143 =>
				ret := to_sfixed(-0.79863551, ret);
			when 144 =>
				ret := to_sfixed(-0.80901699, ret);
			when 145 =>
				ret := to_sfixed(-0.81915204, ret);
			when 146 =>
				ret := to_sfixed(-0.82903757, ret);
			when 147 =>
				ret := to_sfixed(-0.83867057, ret);
			when 148 =>
				ret := to_sfixed(-0.8480481, ret);
			when 149 =>
				ret := to_sfixed(-0.8571673, ret);
			when 150 =>
				ret := to_sfixed(-0.8660254, ret);
			when 151 =>
				ret := to_sfixed(-0.87461971, ret);
			when 152 =>
				ret := to_sfixed(-0.88294759, ret);
			when 153 =>
				ret := to_sfixed(-0.89100652, ret);
			when 154 =>
				ret := to_sfixed(-0.89879405, ret);
			when 155 =>
				ret := to_sfixed(-0.90630779, ret);
			when 156 =>
				ret := to_sfixed(-0.91354546, ret);
			when 157 =>
				ret := to_sfixed(-0.92050485, ret);
			when 158 =>
				ret := to_sfixed(-0.92718385, ret);
			when 159 =>
				ret := to_sfixed(-0.93358043, ret);
			when 160 =>
				ret := to_sfixed(-0.93969262, ret);
			when 161 =>
				ret := to_sfixed(-0.94551858, ret);
			when 162 =>
				ret := to_sfixed(-0.95105652, ret);
			when 163 =>
				ret := to_sfixed(-0.95630476, ret);
			when 164 =>
				ret := to_sfixed(-0.9612617, ret);
			when 165 =>
				ret := to_sfixed(-0.96592583, ret);
			when 166 =>
				ret := to_sfixed(-0.97029573, ret);
			when 167 =>
				ret := to_sfixed(-0.97437006, ret);
			when 168 =>
				ret := to_sfixed(-0.9781476, ret);
			when 169 =>
				ret := to_sfixed(-0.98162718, ret);
			when 170 =>
				ret := to_sfixed(-0.98480775, ret);
			when 171 =>
				ret := to_sfixed(-0.98768834, ret);
			when 172 =>
				ret := to_sfixed(-0.99026807, ret);
			when 173 =>
				ret := to_sfixed(-0.99254615, ret);
			when 174 =>
				ret := to_sfixed(-0.9945219, ret);
			when 175 =>
				ret := to_sfixed(-0.9961947, ret);
			when 176 =>
				ret := to_sfixed(-0.99756405, ret);
			when 177 =>
				ret := to_sfixed(-0.99862953, ret);
			when 178 =>
				ret := to_sfixed(-0.99939083, ret);
			when 179 =>
				ret := to_sfixed(-0.9998477, ret);
			when others =>
				ret := to_sfixed(0.0, ret);
		end case;
		return ret; 
	end cos;
end package;